module sirv_gnrl_ram #(
    parameter DP = 32,
    parameter DW = 32,
    parameter FORCE_X2ZERO = 1,
    parameter MW = 4,
    parameter AW = 15
) (
    
)